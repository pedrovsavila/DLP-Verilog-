module n_b (input [3:0] b,
			  output [3:0] out
			 );
			 
		assign out = ~b;
	
endmodule
				
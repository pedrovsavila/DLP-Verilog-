module myAND ( input A,B,
					output X  );

assign X = A & B;
					
endmodule

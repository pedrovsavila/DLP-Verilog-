module mySUM (
					input signed [3:0] A, B,
					output signed [4:0] X
					);
assign X = A + B;


endmodule
